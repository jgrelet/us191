netcdf test-dboceano-tsg {
dimensions:
	TIME = 5 ;
	LEVEL = 1 ;
	LATITUDE = 5 ;
	LONGITUDE = 5 ;
	POSITION = 5 ;
	STRING256 = 256 ;
	STRING14 = 14 ;
	STRING8 = 8 ;
	STRING4 = 4 ;
	N1 = 1 ;
variables:
	char REFERENCE_DATE_TIME(STRING14) ;
		REFERENCE_DATE_TIME:long_name = "ORIGIN OF TIME" ;
		REFERENCE_DATE_TIME:conventions = "yyyymmddHHMMSS" ;
		REFERENCE_DATE_TIME:comment = "Reference date for julian days origin" ;
	char DATE(TIME, STRING14) ;
		DATE:long_name = "DATE OF MAINS INSTRUMENT MEASUREMENT" ;
		DATE:conventions = "yyyymmddHHMMSS" ;
		DATE:axis = "T" ;
		DATE:comment = "This is the original data describing the date, it must not be lost" ;
		DATE:coordinate = "TIME" ;
	double TIME(TIME) ;
		TIME:long_name = "DECIMAL JULIAN DAY (UTC) OF EACH MEASUREMENT" ;
		TIME:standard_name = "time" ;
		TIME:units = "days since 1950-01-01T00:00:00Z" ;
		TIME:conventions = "Relative julian days with decimal part (as parts of the day) from REFERENCE_DATE_TIME" ;
		TIME:valid_min = 0. ;
		TIME:valid_max = 90000. ;
		TIME:format = "%9.5lf" ;
		TIME:epic_code = 601. ;
		TIME:axis = "T" ;
		TIME:comment = "Julian day of the measurement" ;
		TIME:coordinate = "TIME" ;
	byte TIME_QC(TIME) ;
		TIME_QC:long_name = "QUALITY FLAG OF TIME" ;
		TIME_QC:conventions = "OceanSITES reference table 2" ;
		TIME_QC:valid_min = 0b ;
		TIME_QC:valid_max = 9b ;
		TIME_QC:format = "%1d" ;
		TIME_QC:comment = "Quality flag for each TIME value." ;
		TIME_QC:default_value = 0b ;
		TIME_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		TIME_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float LATITUDE(LATITUDE) ;
		LATITUDE:long_name = "LATITUDE OF THE MEASUREMENT" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degree_north" ;
		LATITUDE:valid_min = -90.f ;
		LATITUDE:valid_max = 90.f ;
		LATITUDE:format = "%+8.4lf" ;
		LATITUDE:_FillValue = 99999.f ;
		LATITUDE:epic_code = 500.f ;
		LATITUDE:axis = "Y" ;
		LATITUDE:comment = "Latitude of the measurement (decimal)" ;
		LATITUDE:coordinate = "LATITUDE" ;
	float LONGITUDE(LONGITUDE) ;
		LONGITUDE:long_name = "LONGITUDE OF THE MEASUREMENT" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degree_east" ;
		LONGITUDE:valid_min = -180.f ;
		LONGITUDE:valid_max = 180.f ;
		LONGITUDE:format = "%+9.4lf" ;
		LONGITUDE:_FillValue = 99999.f ;
		LONGITUDE:epic_code = 501.f ;
		LONGITUDE:axis = "X" ;
		LONGITUDE:comment = "Longitude of the measurement (decimal)" ;
		LONGITUDE:coordinate = "LONGITUDE" ;
	byte POSITION_QC(POSITION) ;
		POSITION_QC:long_name = "QUALITY FLAG OF POSITION" ;
		POSITION_QC:conventions = "OceanSITES reference table 2" ;
		POSITION_QC:valid_min = 0b ;
		POSITION_QC:valid_max = 9b ;
		POSITION_QC:format = "%1d" ;
		POSITION_QC:comment = "Quality flag for each LATITUDE and LONGITUDE value." ;
		POSITION_QC:default_value = 0b ;
		POSITION_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		POSITION_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float SSJT(TIME, LEVEL) ;
		SSJT:long_name = "SEA SURFACE WATER JACKET TEMPERATURE" ;
		SSJT:standard_name = "sea_water_temperature" ;
		SSJT:units = "degree_Celsius" ;
		SSJT:valid_min = -1.5f ;
		SSJT:valid_max = 38.f ;
		SSJT:format = "%6.3lf" ;
		SSJT:_FillValue = 99999.f ;
		SSJT:resolution = 0.001f ;
		SSJT:comment = "Ocean temperature" ;
		SSJT:coordinate = "TIME" ;
	byte SSJT_QC(TIME, LEVEL) ;
		SSJT_QC:long_name = "QUALITY FLAG" ;
		SSJT_QC:conventions = "OceanSITES reference table 2" ;
		SSJT_QC:valid_min = 0b ;
		SSJT_QC:valid_max = 9b ;
		SSJT_QC:format = "%1d" ;
		SSJT_QC:comment = "Quality flag for each Ocean temperature value" ;
		SSJT_QC:default_value = 0b ;
		SSJT_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSJT_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float SSJT_CAL(TIME, LEVEL) ;
		SSJT_CAL:long_name = "SEA SURFACE WATER JACKET TEMPERATURE CALIBRATED" ;
		SSJT_CAL:standard_name = "sea_water_temperature" ;
		SSJT_CAL:units = "degree_Celsius" ;
		SSJT_CAL:valid_min = 99999.f ;
		SSJT_CAL:valid_max = 99999.f ;
		SSJT_CAL:format = "%6.3lf" ;
		SSJT_CAL:_FillValue = 99999.f ;
		SSJT_CAL:comment = "Ocean temperature calibrated" ;
	float SSJT_ADJUSTED(TIME, LEVEL) ;
		SSJT_ADJUSTED:long_name = "SEA SURFACE WATER JACKET TEMPERATURE ADJUSTED" ;
		SSJT_ADJUSTED:standard_name = "sea_water_temperature" ;
		SSJT_ADJUSTED:units = "degree_Celsius" ;
		SSJT_ADJUSTED:valid_min = 99999.f ;
		SSJT_ADJUSTED:valid_max = 99999.f ;
		SSJT_ADJUSTED:format = "%6.3lf" ;
		SSJT_ADJUSTED:_FillValue = 99999.f ;
		SSJT_ADJUSTED:comment = "Adjusted Ocean temperature" ;
	float SSJT_ADJUSTED_ERROR(TIME, LEVEL) ;
		SSJT_ADJUSTED_ERROR:long_name = "ERROR ON SEA SURFACE WATER JACKET TEMPERATURE ADJUSTED" ;
		SSJT_ADJUSTED_ERROR:standard_name = "sea_water_temperature" ;
		SSJT_ADJUSTED_ERROR:units = "degree_Celsius" ;
		SSJT_ADJUSTED_ERROR:valid_min = 99999.f ;
		SSJT_ADJUSTED_ERROR:valid_max = 99999.f ;
		SSJT_ADJUSTED_ERROR:format = "%6.3lf" ;
		SSJT_ADJUSTED_ERROR:_FillValue = 99999.f ;
		SSJT_ADJUSTED_ERROR:comment = "Error on adjusted Ocean temperature" ;
	byte SSJT_ADJUSTED_QC(TIME, LEVEL) ;
		SSJT_ADJUSTED_QC:long_name = "QUALITY FLAG" ;
		SSJT_ADJUSTED_QC:conventions = "OceanSITES reference table 2" ;
		SSJT_ADJUSTED_QC:valid_min = 0b ;
		SSJT_ADJUSTED_QC:valid_max = 9b ;
		SSJT_ADJUSTED_QC:format = "%1d" ;
		SSJT_ADJUSTED_QC:comment = "Quality flag applied on adjusted Ocean temperature" ;
		SSJT_ADJUSTED_QC:default_value = 0b ;
		SSJT_ADJUSTED_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSJT_ADJUSTED_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	char SSJT_ADJUSTED_HIST(STRING256) ;
		SSJT_ADJUSTED_HIST:long_name = "ADJUSTED SEA SURFACE WATER JACKET TEMPERATURE PROCESSING HISTORY" ;
		SSJT_ADJUSTED_HIST:comment = "Adjusted Ocean temperature processing history" ;
	float SSTP(TIME, LEVEL) ;
		SSTP:long_name = "SEA SURFACE WATER TEMPERATURE" ;
		SSTP:standard_name = "sea_water_temperature" ;
		SSTP:units = "degree_Celsius" ;
		SSTP:valid_min = -1.5f ;
		SSTP:valid_max = 38.f ;
		SSTP:format = "%6.3lf" ;
		SSTP:_FillValue = 99999.f ;
		SSTP:resolution = 0.001f ;
		SSTP:comment = "Sea surface Ocean temperature" ;
		SSTP:coordinate = "TIME" ;
	byte SSTP_QC(TIME, LEVEL) ;
		SSTP_QC:long_name = "QUALITY FLAG" ;
		SSTP_QC:conventions = "OceanSITES reference table 2" ;
		SSTP_QC:valid_min = 0b ;
		SSTP_QC:valid_max = 9b ;
		SSTP_QC:format = "%1d" ;
		SSTP_QC:comment = "Quality flag for each Sea surface Ocean temperature value" ;
		SSTP_QC:default_value = 0b ;
		SSTP_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSTP_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float SSTP_CAL(TIME, LEVEL) ;
		SSTP_CAL:long_name = "SEA SURFACE WATER TEMPERATURE CALIBRATED" ;
		SSTP_CAL:standard_name = "sea_water_temperature" ;
		SSTP_CAL:units = "degree_Celsius" ;
		SSTP_CAL:valid_min = 99999.f ;
		SSTP_CAL:valid_max = 99999.f ;
		SSTP_CAL:format = "%6.3lf" ;
		SSTP_CAL:_FillValue = 99999.f ;
		SSTP_CAL:comment = "Sea surface Ocean temperature calibrated" ;
	float SSTP_ADJUSTED(TIME, LEVEL) ;
		SSTP_ADJUSTED:long_name = "SEA SURFACE WATER TEMPERATURE ADJUSTED" ;
		SSTP_ADJUSTED:standard_name = "sea_water_temperature" ;
		SSTP_ADJUSTED:units = "degree_Celsius" ;
		SSTP_ADJUSTED:valid_min = 99999.f ;
		SSTP_ADJUSTED:valid_max = 99999.f ;
		SSTP_ADJUSTED:format = "%6.3lf" ;
		SSTP_ADJUSTED:_FillValue = 99999.f ;
		SSTP_ADJUSTED:comment = "Adjusted Sea surface Ocean temperature" ;
	float SSTP_ADJUSTED_ERROR(TIME, LEVEL) ;
		SSTP_ADJUSTED_ERROR:long_name = "ERROR ON SEA SURFACE WATER TEMPERATURE ADJUSTED" ;
		SSTP_ADJUSTED_ERROR:standard_name = "sea_water_temperature" ;
		SSTP_ADJUSTED_ERROR:units = "degree_Celsius" ;
		SSTP_ADJUSTED_ERROR:valid_min = 99999.f ;
		SSTP_ADJUSTED_ERROR:valid_max = 99999.f ;
		SSTP_ADJUSTED_ERROR:format = "%6.3lf" ;
		SSTP_ADJUSTED_ERROR:_FillValue = 99999.f ;
		SSTP_ADJUSTED_ERROR:comment = "Error on adjusted Sea surface Ocean temperature" ;
	byte SSTP_ADJUSTED_QC(TIME, LEVEL) ;
		SSTP_ADJUSTED_QC:long_name = "QUALITY FLAG" ;
		SSTP_ADJUSTED_QC:conventions = "OceanSITES reference table 2" ;
		SSTP_ADJUSTED_QC:valid_min = 0b ;
		SSTP_ADJUSTED_QC:valid_max = 9b ;
		SSTP_ADJUSTED_QC:format = "%1d" ;
		SSTP_ADJUSTED_QC:comment = "Quality flag applied on adjusted Sea surface Ocean temperature" ;
		SSTP_ADJUSTED_QC:default_value = 0b ;
		SSTP_ADJUSTED_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSTP_ADJUSTED_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	char SSTP_ADJUSTED_HIST(STRING256) ;
		SSTP_ADJUSTED_HIST:long_name = "ADJUSTED SEA SURFACE WATER TEMPERATURE PROCESSING HISTORY" ;
		SSTP_ADJUSTED_HIST:comment = "Adjusted Sea surface Ocean temperature processing history" ;
	float SSPS(TIME, LEVEL) ;
		SSPS:long_name = "SEA SURFACE PRACTICAL SALINITY" ;
		SSPS:standard_name = "sea_water_salinity" ;
		SSPS:units = "psu" ;
		SSPS:valid_min = -1.5f ;
		SSPS:valid_max = 38.f ;
		SSPS:format = "%6.3lf" ;
		SSPS:_FillValue = 99999.f ;
		SSPS:resolution = 0.001f ;
		SSPS:comment = "Ocean salinity" ;
		SSPS:coordinate = "TIME" ;
	byte SSPS_QC(TIME, LEVEL) ;
		SSPS_QC:long_name = "QUALITY FLAG" ;
		SSPS_QC:conventions = "OceanSITES reference table 2" ;
		SSPS_QC:valid_min = 0b ;
		SSPS_QC:valid_max = 9b ;
		SSPS_QC:format = "%1d" ;
		SSPS_QC:comment = "Quality flag for each Ocean salinity value" ;
		SSPS_QC:default_value = 0b ;
		SSPS_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSPS_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float SSPS_CAL(TIME, LEVEL) ;
		SSPS_CAL:long_name = "SEA SURFACE PRACTICAL SALINITY CALIBRATED" ;
		SSPS_CAL:standard_name = "sea_water_salinity" ;
		SSPS_CAL:units = "psu" ;
		SSPS_CAL:valid_min = 99999.f ;
		SSPS_CAL:valid_max = 99999.f ;
		SSPS_CAL:format = "%6.3lf" ;
		SSPS_CAL:_FillValue = 99999.f ;
		SSPS_CAL:comment = "Ocean salinity calibrated" ;
	float SSPS_ADJUSTED(TIME, LEVEL) ;
		SSPS_ADJUSTED:long_name = "SEA SURFACE PRACTICAL SALINITY ADJUSTED" ;
		SSPS_ADJUSTED:standard_name = "sea_water_salinity" ;
		SSPS_ADJUSTED:units = "psu" ;
		SSPS_ADJUSTED:valid_min = 99999.f ;
		SSPS_ADJUSTED:valid_max = 99999.f ;
		SSPS_ADJUSTED:format = "%6.3lf" ;
		SSPS_ADJUSTED:_FillValue = 99999.f ;
		SSPS_ADJUSTED:comment = "Adjusted Ocean salinity" ;
	float SSPS_ADJUSTED_ERROR(TIME, LEVEL) ;
		SSPS_ADJUSTED_ERROR:long_name = "ERROR ON SEA SURFACE PRACTICAL SALINITY ADJUSTED" ;
		SSPS_ADJUSTED_ERROR:standard_name = "sea_water_salinity" ;
		SSPS_ADJUSTED_ERROR:units = "psu" ;
		SSPS_ADJUSTED_ERROR:valid_min = 99999.f ;
		SSPS_ADJUSTED_ERROR:valid_max = 99999.f ;
		SSPS_ADJUSTED_ERROR:format = "%6.3lf" ;
		SSPS_ADJUSTED_ERROR:_FillValue = 99999.f ;
		SSPS_ADJUSTED_ERROR:comment = "Error on adjusted Ocean salinity" ;
	byte SSPS_ADJUSTED_QC(TIME, LEVEL) ;
		SSPS_ADJUSTED_QC:long_name = "QUALITY FLAG" ;
		SSPS_ADJUSTED_QC:conventions = "OceanSITES reference table 2" ;
		SSPS_ADJUSTED_QC:valid_min = 0b ;
		SSPS_ADJUSTED_QC:valid_max = 9b ;
		SSPS_ADJUSTED_QC:format = "%1d" ;
		SSPS_ADJUSTED_QC:comment = "Quality flag applied on adjusted Ocean salinity" ;
		SSPS_ADJUSTED_QC:default_value = 0b ;
		SSPS_ADJUSTED_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		SSPS_ADJUSTED_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	char SSPS_ADJUSTED_HIST(STRING256) ;
		SSPS_ADJUSTED_HIST:long_name = "ADJUSTED SEA SURFACE PRACTICAL SALINITY PROCESSING HISTORY" ;
		SSPS_ADJUSTED_HIST:comment = "Adjusted Ocean salinity processing history" ;
	float PRES(TIME, LEVEL) ;
		PRES:long_name = "SEA WATER PRESSURE" ;
		PRES:standard_name = "sea water pressure" ;
		PRES:units = "decibard" ;
		PRES:positive = "down" ;
		PRES:format = "%7.2lf" ;
		PRES:_FillValue = 99999.f ;
		PRES:axis = "Z" ;
		PRES:comment = "Pressure of the measurement" ;
		PRES:coordinate = "LEVEL" ;
	byte PRES_QC(TIME, LEVEL) ;
		PRES_QC:long_name = "QUALITY FLAG" ;
		PRES_QC:conventions = "OceanSITES reference table 2" ;
		PRES_QC:valid_min = 0b ;
		PRES_QC:valid_max = 9b ;
		PRES_QC:format = "%1d" ;
		PRES_QC:comment = "Quality flag for each level value" ;
		PRES_QC:default_value = 0b ;
		PRES_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		PRES_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;
	float DEPH(TIME, LEVEL) ;
		DEPH:long_name = "SEA WATER DEPH" ;
		DEPH:standard_name = "deph" ;
		DEPH:units = "m" ;
		DEPH:positive = "up" ;
		DEPH:format = "%7.2lf" ;
		DEPH:_FillValue = 99999.f ;
		DEPH:axis = "Z" ;
		DEPH:comment = "Deph of the measurement" ;
		DEPH:coordinate = "LEVEL" ;
	byte DEPH_QC(TIME, LEVEL) ;
		DEPH_QC:long_name = "QUALITY FLAG" ;
		DEPH_QC:conventions = "OceanSITES reference table 2" ;
		DEPH_QC:valid_min = 0b ;
		DEPH_QC:valid_max = 9b ;
		DEPH_QC:format = "%1d" ;
		DEPH_QC:comment = "Quality flag for each level value" ;
		DEPH_QC:default_value = 0b ;
		DEPH_QC:flag_values = "0, 1, 2, 3, 4, 5, 7, 8, 9" ;
		DEPH_QC:flag_meanings = "no_qc_performed, good_data, probably_good_data, bad_data_that_are_potentially_correctable, bad_data, value_changed, not_used, nominal_value, interpolated_value, missing_value" ;

// global attributes:
		:cycle_mesure = "TOUCAN-TEST" ;
		:platform_name = "TOUCAN" ;
		:call_sign = "FNAV" ;
		:wmo_platform_code = "35A9" ;
		:project_name = "ORE-SSS" ;
		:platform_code = "FNAV" ;
		:type_instrument = "SBE21" ;
		:type_position = "GPS" ;
		:number_instrument = "3196" ;
		:data_type = "trajectory" ;
		:data_mode = "N/A" ;
		:time_coverage_start = "2007-07-18T08:40:00Z" ;
		:time_coverage_end = "2007-09-07T09:10:00Z" ;
		:netcdf_version = "3.6" ;
		:conventions = "OceanSITES 1.1, CF1.4" ;
		:date_update = "2010-06-09T15:55:34Z" ;
		:data_restrictions = "N/A" ;
		:pi_name = "Thierry Delcroix" ;
		:author = "Jacques Grelet" ;
		:data_assembly_center = "N/A" ;
		:processing_state = "2C+" ;
		:comment = "N/A" ;
data:

 REFERENCE_DATE_TIME = "19500101000000" ;

 DATE =
  "00570813034500",
  "00570813035000",
  "00570813035500",
  "00570813040000",
  "00570813040500" ;

 TIME = 21045.15625, 21045.1597222222, 21045.1631944445, 21045.1666666666, 
    21045.1701388889 ;

 TIME_QC = -127, -127, -127, -127, -127 ;

 LATITUDE = 16.90657, 16.89335, 16.88023, 16.86723, 16.85425 ;

 LONGITUDE = -64.14038, -64.12425, -64.10775, -64.09133, -64.07475 ;

 POSITION_QC = -127, -127, -127, -127, -127 ;

 SSJT =
  29.185,
  29.241,
  29.252,
  29.266,
  29.261 ;

 SSJT_QC =
  0,
  0,
  0,
  0,
  0 ;

 SSJT_CAL =
  _,
  _,
  _,
  _,
  _ ;

 SSJT_ADJUSTED =
  _,
  _,
  _,
  _,
  _ ;

 SSJT_ADJUSTED_ERROR =
  _,
  _,
  _,
  _,
  _ ;

 SSJT_ADJUSTED_QC =
  0,
  0,
  0,
  0,
  0 ;

 SSJT_ADJUSTED_HIST = "" ;

 SSTP =
  29.085,
  29.141,
  29.152,
  29.166,
  29.161 ;

 SSTP_QC =
  1,
  1,
  1,
  1,
  1 ;

 SSTP_CAL =
  29.086,
  29.142,
  29.153,
  29.267,
  29.162 ;

 SSTP_ADJUSTED =
  29.087,
  29.143,
  29.153,
  29.268,
  29.163 ;

 SSTP_ADJUSTED_ERROR =
  _,
  _,
  _,
  _,
  _ ;

 SSTP_ADJUSTED_QC =
  5,
  5,
  5,
  5,
  5 ;

 SSTP_ADJUSTED_HIST = "" ;

 SSPS =
  35.168,
  35.173,
  35.142,
  35.095,
  35.073 ;

 SSPS_QC =
  1,
  1,
  1,
  1,
  1 ;

 SSPS_CAL =
  35.169,
  35.174,
  35.143,
  35.096,
  35.074 ;

 SSPS_ADJUSTED =
  35.17,
  35.175,
  35.143,
  35.097,
  35.075 ;

 SSPS_ADJUSTED_ERROR =
  _,
  _,
  _,
  _,
  _ ;

 SSPS_ADJUSTED_QC =
  5,
  5,
  5,
  5,
  5 ;

 SSPS_ADJUSTED_HIST = "" ;

 PRES =
  _,
  _,
  _,
  _,
  _ ;

 PRES_QC =
  -127,
  -127,
  -127,
  -127,
  -127 ;

 DEPH =
  _,
  _,
  _,
  _,
  _ ;

 DEPH_QC =
  -127,
  -127,
  -127,
  -127,
  -127 ;
}
