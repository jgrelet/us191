netcdf us191 {
dimensions:
	x = 4 ;
	y = 6 ;
	level = 2 ;
	latitude = 6 ;
	longitude = 12 ;	
        time = UNLIMITED ; // (2 currently)
variables:
	double x(x, y) ;
		x:test_double_att = 3.14159 ;
		x:test_float_att = 3.1416f ;
		x:test_int_att = 3 ;
		x:test_short_att = 5s, 7s ;
		x:test_uchar_att = 100b ;
		x:test_schar_att = -100b ;
		x:test_text_att = "abcdefghijklmnopqrstuvwxyz" ;
		x:new_att = "0" ;
	double test_singleton ;		
	double test_1D(y) ;
      	double test_2D(x, y) ;
		test_2D:_FillValue = -1. ;
		test_2D:missing_value = -1. ;
	short temp(x, y) ;
		temp:scale_factor = 1.8 ;
		temp:add_offset = 32. ;
	float test_2D_float(x, y) ;
	double test_var3(x) ;
	float a(x, y) ;
		a:missing_value = 9999.f ;
	float b(x, y) ;
		b:_FillValue = 9999.f ;
	int test_2D_int ;
		test_2D_int:_FillValue = -1 ;
	short test_2D_short ;
	double time(time) ;
		time:long_name = "Time since initial condition" ;
		time:units = "days since 1950-01-01T00:00:00Z" ;
		time:cartesian_axis = "T" ;
	float latitude(latitude) ;
		latitude:units = "degrees_north" ;
	float longitude(longitude) ;
		longitude:units = "degrees_east" ;
	float pressure(time, level, latitude, longitude) ;
		pressure:units = "hPa" ;
	float temperature(time, level, latitude, longitude) ;
		temperature:units = "celsius" ;
		temperature:missing_value = 32000 ;  // of type short //
		temperature:long_name = "SEA SURFACE TEMPERATURE" ;
		temperature:add_offset = 10.0f ;
		temperature:scale_factor = 2.f ; 
	//temperature:add_offset = 20.0f ;//  
	//	temperature:scale_factor = .0005f ;// 

// global attributes:
		:test_double_att = 3.14159 ;
		:history = "24-Dec-2011 19:30:41" ;
		:date = "12242011T193041Z" ;

data:

 x =
  _ ;

 test_singleton = 3.14159 ;

 test_1D = 1.1, 1.2, 1.3, 1.4, 1.5, 1.6 ;

 test_2D =
  0.1, 0.2, 0.3, 0.4, 0.5, 0.6, 
  0.7, 0.8, 0.9, 1, 1.1, 1.2, 
  1.3, 1.4, 1.5, 1.6, 1.7, 1.8, 
  1.9, 2, 2.1, 2.2, 2.3, 2.4 ;

 time = 47449.9583333333, 47450.9583333333 ;

 latitude = 25, 30, 35, 40, 45, 50 ;

 longitude = -125, -120, -115, -110, -105, -100, -95, -90, -85, -80, -75, -70 ;

 pressure =
  900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911,
  912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923,
  924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935,
  936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947,
  948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959,
  960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971,
  972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983,
  984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995,
  996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007,
  1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019,
  1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031,
  1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043,
  900, 901, 902, 903, 904, 905, 906, 907, 908, 909, 910, 911,
  912, 913, 914, 915, 916, 917, 918, 919, 920, 921, 922, 923,
  924, 925, 926, 927, 928, 929, 930, 931, 932, 933, 934, 935,
  936, 937, 938, 939, 940, 941, 942, 943, 944, 945, 946, 947,
  948, 949, 950, 951, 952, 953, 954, 955, 956, 957, 958, 959,
  960, 961, 962, 963, 964, 965, 966, 967, 968, 969, 970, 971,
  972, 973, 974, 975, 976, 977, 978, 979, 980, 981, 982, 983,
  984, 985, 986, 987, 988, 989, 990, 991, 992, 993, 994, 995,
  996, 997, 998, 999, 1000, 1001, 1002, 1003, 1004, 1005, 1006, 1007,
  1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1018, 1019,
  1020, 1021, 1022, 1023, 1024, 1025, 1026, 1027, 1028, 1029, 1030, 1031,
  1032, 1033, 1034, 1035, 1036, 1037, 1038, 1039, 1040, 1041, 1042, 1043 ;

 temperature =
  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20,
  21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32,
  33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44,
  45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56,
  57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68,
  69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80,
  81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92,
  93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104,
  105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116,
  117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128,
  129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140,
  141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152,
  9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20,
  21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32,
  33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44,
  45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56,
  57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68,
  69, 70, 71, 72, 73, 74, 75, 76, 77, 78, 79, 80,
  81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92,
  93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104,
  105, 106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116,
  117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128,
  129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140,
  141, 142, 143, 144, 145, 146, 147, 148, 149, 150, 151, 152 ;

}
